module weight_rom (
    input clk,
    input reset,
    output reg [15:0] data_out_0,
    output reg [15:0] data_out_1,
    output reg [15:0] data_out_2,
    output reg [15:0] data_out_3,
    output reg [15:0] data_out_4,
    output reg [15:0] data_out_5,
    output reg [15:0] data_out_6,
    output reg [15:0] data_out_7,
    output reg [15:0] data_out_8,
    output reg [15:0] data_out_9,
    output reg [15:0] data_out_10,
    output reg [15:0] data_out_11,
    output reg [15:0] data_out_12,
    output reg [15:0] data_out_13,
    output reg [15:0] data_out_14,
    output reg [15:0] data_out_15,
    output reg [15:0] data_out_16,
    output reg [15:0] data_out_17,
    output reg [15:0] data_out_18,
    output reg [15:0] data_out_19,
    output reg [15:0] data_out_20,
    output reg [15:0] data_out_21,
    output reg [15:0] data_out_22,
    output reg [15:0] data_out_23,
    output reg [15:0] data_out_24,
    output reg [15:0] data_out_25,
    output reg [15:0] data_out_26,
    output reg [15:0] data_out_27,
    output reg [15:0] data_out_28,
    output reg [15:0] data_out_29,
    output reg [15:0] data_out_30,
    output reg [15:0] data_out_31,
    output reg [15:0] data_out_32,
    output reg [15:0] data_out_33,
    output reg [15:0] data_out_34,
    output reg [15:0] data_out_35,
    output reg [15:0] data_out_36,
    output reg [15:0] data_out_37,
    output reg [15:0] data_out_38,
    output reg [15:0] data_out_39,
    output reg [15:0] data_out_40,
    output reg [15:0] data_out_41,
    output reg [15:0] data_out_42,
    output reg [15:0] data_out_43,
    output reg [15:0] data_out_44,
    output reg [15:0] data_out_45,
    output reg [15:0] data_out_46,
    output reg [15:0] data_out_47,
    output reg [15:0] data_out_48,
    output reg [15:0] data_out_49,
    output reg [15:0] data_out_50,
    output reg [15:0] data_out_51,
    output reg [15:0] data_out_52,
    output reg [15:0] data_out_53,
    output reg [15:0] data_out_54,
    output reg [15:0] data_out_55,
    output reg [15:0] data_out_56,
    output reg [15:0] data_out_57,
    output reg [15:0] data_out_58,
    output reg [15:0] data_out_59,
    output reg [15:0] data_out_60,
    output reg [15:0] data_out_61,
    output reg [15:0] data_out_62,
    output reg [15:0] data_out_63,
    output reg [15:0] data_out_64,
    output reg [15:0] data_out_65,
    output reg [15:0] data_out_66,
    output reg [15:0] data_out_67,
    output reg [15:0] data_out_68,
    output reg [15:0] data_out_69,
    output reg [15:0] data_out_70,
    output reg [15:0] data_out_71,
    output reg [15:0] data_out_72,
    output reg [15:0] data_out_73,
    output reg [15:0] data_out_74,
    output reg [15:0] data_out_75,
    output reg [15:0] data_out_76,
    output reg [15:0] data_out_77,
    output reg [15:0] data_out_78,
    output reg [15:0] data_out_79,
    output reg [15:0] data_out_80,
    output reg [15:0] data_out_81,
    output reg [15:0] data_out_82,
    output reg [15:0] data_out_83,
    output reg [15:0] data_out_84,
    output reg [15:0] data_out_85,
    output reg [15:0] data_out_86,
    output reg [15:0] data_out_87,
    output reg [15:0] data_out_88,
    output reg [15:0] data_out_89,
    output reg [15:0] data_out_90,
    output reg [15:0] data_out_91,
    output reg [15:0] data_out_92,
    output reg [15:0] data_out_93,
    output reg [15:0] data_out_94,
    output reg [15:0] data_out_95,
    output reg [15:0] data_out_96,
    output reg [15:0] data_out_97,
    output reg [15:0] data_out_98,
    output reg [15:0] data_out_99,
    output reg [15:0] data_out_100,
    output reg [15:0] data_out_101,
    output reg [15:0] data_out_102,
    output reg [15:0] data_out_103,
    output reg [15:0] data_out_104,
    output reg [15:0] data_out_105,
    output reg [15:0] data_out_106,
    output reg [15:0] data_out_107,
    output reg [15:0] data_out_108,
    output reg [15:0] data_out_109,
    output reg [15:0] data_out_110,
    output reg [15:0] data_out_111,
    output reg [15:0] data_out_112,
    output reg [15:0] data_out_113,
    output reg [15:0] data_out_114,
    output reg [15:0] data_out_115,
    output reg [15:0] data_out_116,
    output reg [15:0] data_out_117,
    output reg [15:0] data_out_118,
    output reg [15:0] data_out_119,
    output reg [15:0] data_out_120,
    output reg [15:0] data_out_121,
    output reg [15:0] data_out_122,
    output reg [15:0] data_out_123,
    output reg [15:0] data_out_124,
    output reg [15:0] data_out_125,
    output reg [15:0] data_out_126,
    output reg [15:0] data_out_127,
    output reg [15:0] data_out_128,
    output reg [15:0] data_out_129,
    output reg [15:0] data_out_130,
    output reg [15:0] data_out_131,
    output reg [15:0] data_out_132,
    output reg [15:0] data_out_133,
    output reg [15:0] data_out_134,
    output reg [15:0] data_out_135,
    output reg [15:0] data_out_136,
    output reg [15:0] data_out_137,
    output reg [15:0] data_out_138,
    output reg [15:0] data_out_139,
    output reg [15:0] data_out_140,
    output reg [15:0] data_out_141,
    output reg [15:0] data_out_142,
    output reg [15:0] data_out_143,
    output reg [15:0] data_out_144,
    output reg [15:0] data_out_145,
    output reg [15:0] data_out_146,
    output reg [15:0] data_out_147,
    output reg [15:0] data_out_148,
    output reg [15:0] data_out_149,
    output reg [15:0] data_out_150,
    output reg [15:0] data_out_151,
    output reg [15:0] data_out_152,
    output reg [15:0] data_out_153,
    output reg [15:0] data_out_154,
    output reg [15:0] data_out_155,
    output reg [15:0] data_out_156,
    output reg [15:0] data_out_157,
    output reg [15:0] data_out_158,
    output reg [15:0] data_out_159,
    output reg [15:0] data_out_160,
    output reg [15:0] data_out_161,
    output reg [15:0] data_out_162,
    output reg [15:0] data_out_163,
    output reg [15:0] data_out_164,
    output reg [15:0] data_out_165,
    output reg [15:0] data_out_166,
    output reg [15:0] data_out_167,
    output reg [15:0] data_out_168,
    output reg [15:0] data_out_169,
    output reg [15:0] data_out_170,
    output reg [15:0] data_out_171,
    output reg [15:0] data_out_172,
    output reg [15:0] data_out_173,
    output reg [15:0] data_out_174,
    output reg [15:0] data_out_175,
    output reg [15:0] data_out_176,
    output reg [15:0] data_out_177,
    output reg [15:0] data_out_178,
    output reg [15:0] data_out_179,
    output reg [15:0] data_out_180,
    output reg [15:0] data_out_181,
    output reg [15:0] data_out_182,
    output reg [15:0] data_out_183,
    output reg [15:0] data_out_184,
    output reg [15:0] data_out_185,
    output reg [15:0] data_out_186,
    output reg [15:0] data_out_187,
    output reg [15:0] data_out_188,
    output reg [15:0] data_out_189,
    output reg [15:0] data_out_190,
    output reg [15:0] data_out_191
);

    // ROM data initialization (example weights for simplicity)
    // Define a 192 x 16-bit memory array
    (* ram_style = "block" *) reg [15:0] rom_data [0:191]; 
	
	// Preload memory from a file during initialization
    initial begin
        $readmemh("weight_rom.hex", rom_data);     // Load the instruction memory from the hex file
    end

    always @(posedge clk or posedge reset) begin
        if (reset) begin
            // Reset logic if needed
        end else begin
            // Fetch data from ROM based on the address
            data_out_0   <= rom_data[0];
			data_out_1   <= rom_data[1];
			data_out_2   <= rom_data[2];
			data_out_3   <= rom_data[3];
			data_out_4   <= rom_data[4];
			data_out_5   <= rom_data[5];
			data_out_6   <= rom_data[6];
			data_out_7   <= rom_data[7];
			data_out_8   <= rom_data[8];
			data_out_9   <= rom_data[9];
			data_out_10  <= rom_data[10];
			data_out_11  <= rom_data[11];
			data_out_12  <= rom_data[12];
			data_out_13  <= rom_data[13];
			data_out_14  <= rom_data[14];
			data_out_15  <= rom_data[15];
			data_out_16  <= rom_data[16];
			data_out_17  <= rom_data[17];
			data_out_18  <= rom_data[18];
			data_out_19  <= rom_data[19];
			data_out_20  <= rom_data[20];
			data_out_21  <= rom_data[21];
			data_out_22  <= rom_data[22];
			data_out_23  <= rom_data[23];
			data_out_24  <= rom_data[24];
			data_out_25  <= rom_data[25];
			data_out_26  <= rom_data[26];
			data_out_27  <= rom_data[27];
			data_out_28  <= rom_data[28];
			data_out_29  <= rom_data[29];
			data_out_30  <= rom_data[30];
			data_out_31  <= rom_data[31];
			data_out_32  <= rom_data[32];
			data_out_33  <= rom_data[33];
			data_out_34  <= rom_data[34];
			data_out_35  <= rom_data[35];
			data_out_36  <= rom_data[36];
			data_out_37  <= rom_data[37];
			data_out_38  <= rom_data[38];
			data_out_39  <= rom_data[39];
			data_out_40  <= rom_data[40];
			data_out_41  <= rom_data[41];
			data_out_42  <= rom_data[42];
			data_out_43  <= rom_data[43];
			data_out_44  <= rom_data[44];
			data_out_45  <= rom_data[45];
			data_out_46  <= rom_data[46];
			data_out_47  <= rom_data[47];
			data_out_48  <= rom_data[48];
			data_out_49  <= rom_data[49];
			data_out_50  <= rom_data[50];
			data_out_51  <= rom_data[51];
			data_out_52  <= rom_data[52];
			data_out_53  <= rom_data[53];
			data_out_54  <= rom_data[54];
			data_out_55  <= rom_data[55];
			data_out_56  <= rom_data[56];
			data_out_57  <= rom_data[57];
			data_out_58  <= rom_data[58];
			data_out_59  <= rom_data[59];
			data_out_60  <= rom_data[60];
			data_out_61  <= rom_data[61];
			data_out_62  <= rom_data[62];
			data_out_63  <= rom_data[63];
			data_out_64  <= rom_data[64];
			data_out_65  <= rom_data[65];
			data_out_66  <= rom_data[66];
			data_out_67  <= rom_data[67];
			data_out_68  <= rom_data[68];
			data_out_69  <= rom_data[69];
			data_out_70  <= rom_data[70];
			data_out_71  <= rom_data[71];
			data_out_72  <= rom_data[72];
			data_out_73  <= rom_data[73];
			data_out_74  <= rom_data[74];
			data_out_75  <= rom_data[75];
			data_out_76  <= rom_data[76];
			data_out_77  <= rom_data[77];
			data_out_78  <= rom_data[78];
			data_out_79  <= rom_data[79];
			data_out_80  <= rom_data[80];
			data_out_81  <= rom_data[81];
			data_out_82  <= rom_data[82];
			data_out_83  <= rom_data[83];
			data_out_84  <= rom_data[84];
			data_out_85  <= rom_data[85];
			data_out_86  <= rom_data[86];
			data_out_87  <= rom_data[87];
			data_out_88  <= rom_data[88];
			data_out_89  <= rom_data[89];
			data_out_90  <= rom_data[90];
			data_out_91  <= rom_data[91];
			data_out_92  <= rom_data[92];
			data_out_93  <= rom_data[93];
			data_out_94  <= rom_data[94];
			data_out_95  <= rom_data[95];
			data_out_96  <= rom_data[96];
			data_out_97  <= rom_data[97];
			data_out_98  <= rom_data[98];
			data_out_99  <= rom_data[99];
			data_out_100 <= rom_data[100];
			data_out_101 <= rom_data[101];
			data_out_102 <= rom_data[102];
			data_out_103 <= rom_data[103];
			data_out_104 <= rom_data[104];
			data_out_105 <= rom_data[105];
			data_out_106 <= rom_data[106];
			data_out_107 <= rom_data[107];
			data_out_108 <= rom_data[108];
			data_out_109 <= rom_data[109];
			data_out_110 <= rom_data[110];
			data_out_111 <= rom_data[111];
			data_out_112 <= rom_data[112];
			data_out_113 <= rom_data[113];
			data_out_114 <= rom_data[114];
			data_out_115 <= rom_data[115];
			data_out_116 <= rom_data[116];
			data_out_117 <= rom_data[117];
			data_out_118 <= rom_data[118];
			data_out_119 <= rom_data[119];
			data_out_120 <= rom_data[120];
			data_out_121 <= rom_data[121];
			data_out_122 <= rom_data[122];
			data_out_123 <= rom_data[123];
			data_out_124 <= rom_data[124];
			data_out_125 <= rom_data[125];
			data_out_126 <= rom_data[126];
			data_out_127 <= rom_data[127];
			data_out_128 <= rom_data[128];
			data_out_129 <= rom_data[129];
			data_out_130 <= rom_data[130];
			data_out_131 <= rom_data[131];
			data_out_132 <= rom_data[132];
			data_out_133 <= rom_data[133];
			data_out_134 <= rom_data[134];
			data_out_135 <= rom_data[135];
			data_out_136 <= rom_data[136];
			data_out_137 <= rom_data[137];
			data_out_138 <= rom_data[138];
			data_out_139 <= rom_data[139];
			data_out_140 <= rom_data[140];
			data_out_141 <= rom_data[141];
			data_out_142 <= rom_data[142];
			data_out_143 <= rom_data[143];
			data_out_144 <= rom_data[144];
			data_out_145 <= rom_data[145];
			data_out_146 <= rom_data[146];
			data_out_147 <= rom_data[147];
			data_out_148 <= rom_data[148];
			data_out_149 <= rom_data[149];
			data_out_150 <= rom_data[150];
			data_out_151 <= rom_data[151];
			data_out_152 <= rom_data[152];
			data_out_153 <= rom_data[153];
			data_out_154 <= rom_data[154];
			data_out_155 <= rom_data[155];
			data_out_156 <= rom_data[156];
			data_out_157 <= rom_data[157];
			data_out_158 <= rom_data[158];
			data_out_159 <= rom_data[159];
			data_out_160 <= rom_data[160];
			data_out_161 <= rom_data[161];
			data_out_162 <= rom_data[162];
			data_out_163 <= rom_data[163];
			data_out_164 <= rom_data[164];
			data_out_165 <= rom_data[165];
			data_out_166 <= rom_data[166];
			data_out_167 <= rom_data[167];
			data_out_168 <= rom_data[168];
			data_out_169 <= rom_data[169];
			data_out_170 <= rom_data[170];
			data_out_171 <= rom_data[171];
			data_out_172 <= rom_data[172];
			data_out_173 <= rom_data[173];
			data_out_174 <= rom_data[174];
			data_out_175 <= rom_data[175];
			data_out_176 <= rom_data[176];
			data_out_177 <= rom_data[177];
			data_out_178 <= rom_data[178];
			data_out_179 <= rom_data[179];
			data_out_180 <= rom_data[180];
			data_out_181 <= rom_data[181];
			data_out_182 <= rom_data[182];
			data_out_183 <= rom_data[183];
			data_out_184 <= rom_data[184];
			data_out_185 <= rom_data[185];
			data_out_186 <= rom_data[186];
			data_out_187 <= rom_data[187];
			data_out_188 <= rom_data[188];
			data_out_189 <= rom_data[189];
			data_out_190 <= rom_data[190];
			data_out_191 <= rom_data[191];

        end
    end
endmodule
