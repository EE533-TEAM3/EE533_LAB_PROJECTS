module NPU_top(
	input clk, reset
    
);

    wire [15:0] wire_weight_from_rom [739:0];
	
	
	
	wire [15:0] wire_hiddenlayer_neuron_result [9:0];
	
	wire [15:0] wire_ReLu_result [9:0];
	
	wire [15:0] output_layer_neuron [9:0];
	
	wire [15:0] final_inference;
	
	wire [63:0] data_in; // used for testing. Eventually, it will be an input port for netfpga data to go thru.
	
	assign data_in = 64'b0000111000111100001000000011100000001100000011000011100000110000;

	

	//instantiate rom with weights
	weight_rom weight_rom(
		.clk(clk),
		.reset(reset),                               
			.data_out_0  (wire_weight_from_rom[0]),
			.data_out_1  (wire_weight_from_rom[1]),
			.data_out_2  (wire_weight_from_rom[2]),
			.data_out_3  (wire_weight_from_rom[3]),
			.data_out_4  (wire_weight_from_rom[4]),
			.data_out_5  (wire_weight_from_rom[5]),
			.data_out_6  (wire_weight_from_rom[6]),
			.data_out_7  (wire_weight_from_rom[7]),
			.data_out_8  (wire_weight_from_rom[8]),
			.data_out_9  (wire_weight_from_rom[9]),
			.data_out_10  (wire_weight_from_rom[10]),
			.data_out_11  (wire_weight_from_rom[11]),
			.data_out_12  (wire_weight_from_rom[12]),
			.data_out_13  (wire_weight_from_rom[13]),
			.data_out_14  (wire_weight_from_rom[14]),
			.data_out_15  (wire_weight_from_rom[15]),
			.data_out_16  (wire_weight_from_rom[16]),
			.data_out_17  (wire_weight_from_rom[17]),
			.data_out_18  (wire_weight_from_rom[18]),
			.data_out_19  (wire_weight_from_rom[19]),
			.data_out_20  (wire_weight_from_rom[20]),
			.data_out_21  (wire_weight_from_rom[21]),
			.data_out_22  (wire_weight_from_rom[22]),
			.data_out_23  (wire_weight_from_rom[23]),
			.data_out_24  (wire_weight_from_rom[24]),
			.data_out_25  (wire_weight_from_rom[25]),
			.data_out_26  (wire_weight_from_rom[26]),
			.data_out_27  (wire_weight_from_rom[27]),
			.data_out_28  (wire_weight_from_rom[28]),
			.data_out_29  (wire_weight_from_rom[29]),
			.data_out_30  (wire_weight_from_rom[30]),
			.data_out_31  (wire_weight_from_rom[31]),
			.data_out_32  (wire_weight_from_rom[32]),
			.data_out_33  (wire_weight_from_rom[33]),
			.data_out_34  (wire_weight_from_rom[34]),
			.data_out_35  (wire_weight_from_rom[35]),
			.data_out_36  (wire_weight_from_rom[36]),
			.data_out_37  (wire_weight_from_rom[37]),
			.data_out_38  (wire_weight_from_rom[38]),
			.data_out_39  (wire_weight_from_rom[39]),
			.data_out_40  (wire_weight_from_rom[40]),
			.data_out_41  (wire_weight_from_rom[41]),
			.data_out_42  (wire_weight_from_rom[42]),
			.data_out_43  (wire_weight_from_rom[43]),
			.data_out_44  (wire_weight_from_rom[44]),
			.data_out_45  (wire_weight_from_rom[45]),
			.data_out_46  (wire_weight_from_rom[46]),
			.data_out_47  (wire_weight_from_rom[47]),
			.data_out_48  (wire_weight_from_rom[48]),
			.data_out_49  (wire_weight_from_rom[49]),
			.data_out_50  (wire_weight_from_rom[50]),
			.data_out_51  (wire_weight_from_rom[51]),
			.data_out_52  (wire_weight_from_rom[52]),
			.data_out_53  (wire_weight_from_rom[53]),
			.data_out_54  (wire_weight_from_rom[54]),
			.data_out_55  (wire_weight_from_rom[55]),
			.data_out_56  (wire_weight_from_rom[56]),
			.data_out_57  (wire_weight_from_rom[57]),
			.data_out_58  (wire_weight_from_rom[58]),
			.data_out_59  (wire_weight_from_rom[59]),
			.data_out_60  (wire_weight_from_rom[60]),
			.data_out_61  (wire_weight_from_rom[61]),
			.data_out_62  (wire_weight_from_rom[62]),
			.data_out_63  (wire_weight_from_rom[63]),
			.data_out_64  (wire_weight_from_rom[64]),
			.data_out_65  (wire_weight_from_rom[65]),
			.data_out_66  (wire_weight_from_rom[66]),
			.data_out_67  (wire_weight_from_rom[67]),
			.data_out_68  (wire_weight_from_rom[68]),
			.data_out_69  (wire_weight_from_rom[69]),
			.data_out_70  (wire_weight_from_rom[70]),
			.data_out_71  (wire_weight_from_rom[71]),
			.data_out_72  (wire_weight_from_rom[72]),
			.data_out_73  (wire_weight_from_rom[73]),
			.data_out_74  (wire_weight_from_rom[74]),
			.data_out_75  (wire_weight_from_rom[75]),
			.data_out_76  (wire_weight_from_rom[76]),
			.data_out_77  (wire_weight_from_rom[77]),
			.data_out_78  (wire_weight_from_rom[78]),
			.data_out_79  (wire_weight_from_rom[79]),
			.data_out_80  (wire_weight_from_rom[80]),
			.data_out_81  (wire_weight_from_rom[81]),
			.data_out_82  (wire_weight_from_rom[82]),
			.data_out_83  (wire_weight_from_rom[83]),
			.data_out_84  (wire_weight_from_rom[84]),
			.data_out_85  (wire_weight_from_rom[85]),
			.data_out_86  (wire_weight_from_rom[86]),
			.data_out_87  (wire_weight_from_rom[87]),
			.data_out_88  (wire_weight_from_rom[88]),
			.data_out_89  (wire_weight_from_rom[89]),
			.data_out_90  (wire_weight_from_rom[90]),
			.data_out_91  (wire_weight_from_rom[91]),
			.data_out_92  (wire_weight_from_rom[92]),
			.data_out_93  (wire_weight_from_rom[93]),
			.data_out_94  (wire_weight_from_rom[94]),
			.data_out_95  (wire_weight_from_rom[95]),
			.data_out_96  (wire_weight_from_rom[96]),
			.data_out_97  (wire_weight_from_rom[97]),
			.data_out_98  (wire_weight_from_rom[98]),
			.data_out_99  (wire_weight_from_rom[99]),
			.data_out_100  (wire_weight_from_rom[100]),
			.data_out_101  (wire_weight_from_rom[101]),
			.data_out_102  (wire_weight_from_rom[102]),
			.data_out_103  (wire_weight_from_rom[103]),
			.data_out_104  (wire_weight_from_rom[104]),
			.data_out_105  (wire_weight_from_rom[105]),
			.data_out_106  (wire_weight_from_rom[106]),
			.data_out_107  (wire_weight_from_rom[107]),
			.data_out_108  (wire_weight_from_rom[108]),
			.data_out_109  (wire_weight_from_rom[109]),
			.data_out_110  (wire_weight_from_rom[110]),
			.data_out_111  (wire_weight_from_rom[111]),
			.data_out_112  (wire_weight_from_rom[112]),
			.data_out_113  (wire_weight_from_rom[113]),
			.data_out_114  (wire_weight_from_rom[114]),
			.data_out_115  (wire_weight_from_rom[115]),
			.data_out_116  (wire_weight_from_rom[116]),
			.data_out_117  (wire_weight_from_rom[117]),
			.data_out_118  (wire_weight_from_rom[118]),
			.data_out_119  (wire_weight_from_rom[119]),
			.data_out_120  (wire_weight_from_rom[120]),
			.data_out_121  (wire_weight_from_rom[121]),
			.data_out_122  (wire_weight_from_rom[122]),
			.data_out_123  (wire_weight_from_rom[123]),
			.data_out_124  (wire_weight_from_rom[124]),
			.data_out_125  (wire_weight_from_rom[125]),
			.data_out_126  (wire_weight_from_rom[126]),
			.data_out_127  (wire_weight_from_rom[127]),
			.data_out_128  (wire_weight_from_rom[128]),
			.data_out_129  (wire_weight_from_rom[129]),
			.data_out_130  (wire_weight_from_rom[130]),
			.data_out_131  (wire_weight_from_rom[131]),
			.data_out_132  (wire_weight_from_rom[132]),
			.data_out_133  (wire_weight_from_rom[133]),
			.data_out_134  (wire_weight_from_rom[134]),
			.data_out_135  (wire_weight_from_rom[135]),
			.data_out_136  (wire_weight_from_rom[136]),
			.data_out_137  (wire_weight_from_rom[137]),
			.data_out_138  (wire_weight_from_rom[138]),
			.data_out_139  (wire_weight_from_rom[139]),
			.data_out_140  (wire_weight_from_rom[140]),
			.data_out_141  (wire_weight_from_rom[141]),
			.data_out_142  (wire_weight_from_rom[142]),
			.data_out_143  (wire_weight_from_rom[143]),
			.data_out_144  (wire_weight_from_rom[144]),
			.data_out_145  (wire_weight_from_rom[145]),
			.data_out_146  (wire_weight_from_rom[146]),
			.data_out_147  (wire_weight_from_rom[147]),
			.data_out_148  (wire_weight_from_rom[148]),
			.data_out_149  (wire_weight_from_rom[149]),
			.data_out_150  (wire_weight_from_rom[150]),
			.data_out_151  (wire_weight_from_rom[151]),
			.data_out_152  (wire_weight_from_rom[152]),
			.data_out_153  (wire_weight_from_rom[153]),
			.data_out_154  (wire_weight_from_rom[154]),
			.data_out_155  (wire_weight_from_rom[155]),
			.data_out_156  (wire_weight_from_rom[156]),
			.data_out_157  (wire_weight_from_rom[157]),
			.data_out_158  (wire_weight_from_rom[158]),
			.data_out_159  (wire_weight_from_rom[159]),
			.data_out_160  (wire_weight_from_rom[160]),
			.data_out_161  (wire_weight_from_rom[161]),
			.data_out_162  (wire_weight_from_rom[162]),
			.data_out_163  (wire_weight_from_rom[163]),
			.data_out_164  (wire_weight_from_rom[164]),
			.data_out_165  (wire_weight_from_rom[165]),
			.data_out_166  (wire_weight_from_rom[166]),
			.data_out_167  (wire_weight_from_rom[167]),
			.data_out_168  (wire_weight_from_rom[168]),
			.data_out_169  (wire_weight_from_rom[169]),
			.data_out_170  (wire_weight_from_rom[170]),
			.data_out_171  (wire_weight_from_rom[171]),
			.data_out_172  (wire_weight_from_rom[172]),
			.data_out_173  (wire_weight_from_rom[173]),
			.data_out_174  (wire_weight_from_rom[174]),
			.data_out_175  (wire_weight_from_rom[175]),
			.data_out_176  (wire_weight_from_rom[176]),
			.data_out_177  (wire_weight_from_rom[177]),
			.data_out_178  (wire_weight_from_rom[178]),
			.data_out_179  (wire_weight_from_rom[179]),
			.data_out_180  (wire_weight_from_rom[180]),
			.data_out_181  (wire_weight_from_rom[181]),
			.data_out_182  (wire_weight_from_rom[182]),
			.data_out_183  (wire_weight_from_rom[183]),
			.data_out_184  (wire_weight_from_rom[184]),
			.data_out_185  (wire_weight_from_rom[185]),
			.data_out_186  (wire_weight_from_rom[186]),
			.data_out_187  (wire_weight_from_rom[187]),
			.data_out_188  (wire_weight_from_rom[188]),
			.data_out_189  (wire_weight_from_rom[189]),
			.data_out_190  (wire_weight_from_rom[190]),
			.data_out_191  (wire_weight_from_rom[191]),
			.data_out_192  (wire_weight_from_rom[192]),
			.data_out_193  (wire_weight_from_rom[193]),
			.data_out_194  (wire_weight_from_rom[194]),
			.data_out_195  (wire_weight_from_rom[195]),
			.data_out_196  (wire_weight_from_rom[196]),
			.data_out_197  (wire_weight_from_rom[197]),
			.data_out_198  (wire_weight_from_rom[198]),
			.data_out_199  (wire_weight_from_rom[199]),
			.data_out_200  (wire_weight_from_rom[200]),
			.data_out_201  (wire_weight_from_rom[201]),
			.data_out_202  (wire_weight_from_rom[202]),
			.data_out_203  (wire_weight_from_rom[203]),
			.data_out_204  (wire_weight_from_rom[204]),
			.data_out_205  (wire_weight_from_rom[205]),
			.data_out_206  (wire_weight_from_rom[206]),
			.data_out_207  (wire_weight_from_rom[207]),
			.data_out_208  (wire_weight_from_rom[208]),
			.data_out_209  (wire_weight_from_rom[209]),
			.data_out_210  (wire_weight_from_rom[210]),
			.data_out_211  (wire_weight_from_rom[211]),
			.data_out_212  (wire_weight_from_rom[212]),
			.data_out_213  (wire_weight_from_rom[213]),
			.data_out_214  (wire_weight_from_rom[214]),
			.data_out_215  (wire_weight_from_rom[215]),
			.data_out_216  (wire_weight_from_rom[216]),
			.data_out_217  (wire_weight_from_rom[217]),
			.data_out_218  (wire_weight_from_rom[218]),
			.data_out_219  (wire_weight_from_rom[219]),
			.data_out_220  (wire_weight_from_rom[220]),
			.data_out_221  (wire_weight_from_rom[221]),
			.data_out_222  (wire_weight_from_rom[222]),
			.data_out_223  (wire_weight_from_rom[223]),
			.data_out_224  (wire_weight_from_rom[224]),
			.data_out_225  (wire_weight_from_rom[225]),
			.data_out_226  (wire_weight_from_rom[226]),
			.data_out_227  (wire_weight_from_rom[227]),
			.data_out_228  (wire_weight_from_rom[228]),
			.data_out_229  (wire_weight_from_rom[229]),
			.data_out_230  (wire_weight_from_rom[230]),
			.data_out_231  (wire_weight_from_rom[231]),
			.data_out_232  (wire_weight_from_rom[232]),
			.data_out_233  (wire_weight_from_rom[233]),
			.data_out_234  (wire_weight_from_rom[234]),
			.data_out_235  (wire_weight_from_rom[235]),
			.data_out_236  (wire_weight_from_rom[236]),
			.data_out_237  (wire_weight_from_rom[237]),
			.data_out_238  (wire_weight_from_rom[238]),
			.data_out_239  (wire_weight_from_rom[239]),
			.data_out_240  (wire_weight_from_rom[240]),
			.data_out_241  (wire_weight_from_rom[241]),
			.data_out_242  (wire_weight_from_rom[242]),
			.data_out_243  (wire_weight_from_rom[243]),
			.data_out_244  (wire_weight_from_rom[244]),
			.data_out_245  (wire_weight_from_rom[245]),
			.data_out_246  (wire_weight_from_rom[246]),
			.data_out_247  (wire_weight_from_rom[247]),
			.data_out_248  (wire_weight_from_rom[248]),
			.data_out_249  (wire_weight_from_rom[249]),
			.data_out_250  (wire_weight_from_rom[250]),
			.data_out_251  (wire_weight_from_rom[251]),
			.data_out_252  (wire_weight_from_rom[252]),
			.data_out_253  (wire_weight_from_rom[253]),
			.data_out_254  (wire_weight_from_rom[254]),
			.data_out_255  (wire_weight_from_rom[255]),
			.data_out_256  (wire_weight_from_rom[256]),
			.data_out_257  (wire_weight_from_rom[257]),
			.data_out_258  (wire_weight_from_rom[258]),
			.data_out_259  (wire_weight_from_rom[259]),
			.data_out_260  (wire_weight_from_rom[260]),
			.data_out_261  (wire_weight_from_rom[261]),
			.data_out_262  (wire_weight_from_rom[262]),
			.data_out_263  (wire_weight_from_rom[263]),
			.data_out_264  (wire_weight_from_rom[264]),
			.data_out_265  (wire_weight_from_rom[265]),
			.data_out_266  (wire_weight_from_rom[266]),
			.data_out_267  (wire_weight_from_rom[267]),
			.data_out_268  (wire_weight_from_rom[268]),
			.data_out_269  (wire_weight_from_rom[269]),
			.data_out_270  (wire_weight_from_rom[270]),
			.data_out_271  (wire_weight_from_rom[271]),
			.data_out_272  (wire_weight_from_rom[272]),
			.data_out_273  (wire_weight_from_rom[273]),
			.data_out_274  (wire_weight_from_rom[274]),
			.data_out_275  (wire_weight_from_rom[275]),
			.data_out_276  (wire_weight_from_rom[276]),
			.data_out_277  (wire_weight_from_rom[277]),
			.data_out_278  (wire_weight_from_rom[278]),
			.data_out_279  (wire_weight_from_rom[279]),
			.data_out_280  (wire_weight_from_rom[280]),
			.data_out_281  (wire_weight_from_rom[281]),
			.data_out_282  (wire_weight_from_rom[282]),
			.data_out_283  (wire_weight_from_rom[283]),
			.data_out_284  (wire_weight_from_rom[284]),
			.data_out_285  (wire_weight_from_rom[285]),
			.data_out_286  (wire_weight_from_rom[286]),
			.data_out_287  (wire_weight_from_rom[287]),
			.data_out_288  (wire_weight_from_rom[288]),
			.data_out_289  (wire_weight_from_rom[289]),
			.data_out_290  (wire_weight_from_rom[290]),
			.data_out_291  (wire_weight_from_rom[291]),
			.data_out_292  (wire_weight_from_rom[292]),
			.data_out_293  (wire_weight_from_rom[293]),
			.data_out_294  (wire_weight_from_rom[294]),
			.data_out_295  (wire_weight_from_rom[295]),
			.data_out_296  (wire_weight_from_rom[296]),
			.data_out_297  (wire_weight_from_rom[297]),
			.data_out_298  (wire_weight_from_rom[298]),
			.data_out_299  (wire_weight_from_rom[299]),
			.data_out_300  (wire_weight_from_rom[300]),
			.data_out_301  (wire_weight_from_rom[301]),
			.data_out_302  (wire_weight_from_rom[302]),
			.data_out_303  (wire_weight_from_rom[303]),
			.data_out_304  (wire_weight_from_rom[304]),
			.data_out_305  (wire_weight_from_rom[305]),
			.data_out_306  (wire_weight_from_rom[306]),
			.data_out_307  (wire_weight_from_rom[307]),
			.data_out_308  (wire_weight_from_rom[308]),
			.data_out_309  (wire_weight_from_rom[309]),
			.data_out_310  (wire_weight_from_rom[310]),
			.data_out_311  (wire_weight_from_rom[311]),
			.data_out_312  (wire_weight_from_rom[312]),
			.data_out_313  (wire_weight_from_rom[313]),
			.data_out_314  (wire_weight_from_rom[314]),
			.data_out_315  (wire_weight_from_rom[315]),
			.data_out_316  (wire_weight_from_rom[316]),
			.data_out_317  (wire_weight_from_rom[317]),
			.data_out_318  (wire_weight_from_rom[318]),
			.data_out_319  (wire_weight_from_rom[319]),
			.data_out_320  (wire_weight_from_rom[320]),
			.data_out_321  (wire_weight_from_rom[321]),
			.data_out_322  (wire_weight_from_rom[322]),
			.data_out_323  (wire_weight_from_rom[323]),
			.data_out_324  (wire_weight_from_rom[324]),
			.data_out_325  (wire_weight_from_rom[325]),
			.data_out_326  (wire_weight_from_rom[326]),
			.data_out_327  (wire_weight_from_rom[327]),
			.data_out_328  (wire_weight_from_rom[328]),
			.data_out_329  (wire_weight_from_rom[329]),
			.data_out_330  (wire_weight_from_rom[330]),
			.data_out_331  (wire_weight_from_rom[331]),
			.data_out_332  (wire_weight_from_rom[332]),
			.data_out_333  (wire_weight_from_rom[333]),
			.data_out_334  (wire_weight_from_rom[334]),
			.data_out_335  (wire_weight_from_rom[335]),
			.data_out_336  (wire_weight_from_rom[336]),
			.data_out_337  (wire_weight_from_rom[337]),
			.data_out_338  (wire_weight_from_rom[338]),
			.data_out_339  (wire_weight_from_rom[339]),
			.data_out_340  (wire_weight_from_rom[340]),
			.data_out_341  (wire_weight_from_rom[341]),
			.data_out_342  (wire_weight_from_rom[342]),
			.data_out_343  (wire_weight_from_rom[343]),
			.data_out_344  (wire_weight_from_rom[344]),
			.data_out_345  (wire_weight_from_rom[345]),
			.data_out_346  (wire_weight_from_rom[346]),
			.data_out_347  (wire_weight_from_rom[347]),
			.data_out_348  (wire_weight_from_rom[348]),
			.data_out_349  (wire_weight_from_rom[349]),
			.data_out_350  (wire_weight_from_rom[350]),
			.data_out_351  (wire_weight_from_rom[351]),
			.data_out_352  (wire_weight_from_rom[352]),
			.data_out_353  (wire_weight_from_rom[353]),
			.data_out_354  (wire_weight_from_rom[354]),
			.data_out_355  (wire_weight_from_rom[355]),
			.data_out_356  (wire_weight_from_rom[356]),
			.data_out_357  (wire_weight_from_rom[357]),
			.data_out_358  (wire_weight_from_rom[358]),
			.data_out_359  (wire_weight_from_rom[359]),
			.data_out_360  (wire_weight_from_rom[360]),
			.data_out_361  (wire_weight_from_rom[361]),
			.data_out_362  (wire_weight_from_rom[362]),
			.data_out_363  (wire_weight_from_rom[363]),
			.data_out_364  (wire_weight_from_rom[364]),
			.data_out_365  (wire_weight_from_rom[365]),
			.data_out_366  (wire_weight_from_rom[366]),
			.data_out_367  (wire_weight_from_rom[367]),
			.data_out_368  (wire_weight_from_rom[368]),
			.data_out_369  (wire_weight_from_rom[369]),
			.data_out_370  (wire_weight_from_rom[370]),
			.data_out_371  (wire_weight_from_rom[371]),
			.data_out_372  (wire_weight_from_rom[372]),
			.data_out_373  (wire_weight_from_rom[373]),
			.data_out_374  (wire_weight_from_rom[374]),
			.data_out_375  (wire_weight_from_rom[375]),
			.data_out_376  (wire_weight_from_rom[376]),
			.data_out_377  (wire_weight_from_rom[377]),
			.data_out_378  (wire_weight_from_rom[378]),
			.data_out_379  (wire_weight_from_rom[379]),
			.data_out_380  (wire_weight_from_rom[380]),
			.data_out_381  (wire_weight_from_rom[381]),
			.data_out_382  (wire_weight_from_rom[382]),
			.data_out_383  (wire_weight_from_rom[383]),
			.data_out_384  (wire_weight_from_rom[384]),
			.data_out_385  (wire_weight_from_rom[385]),
			.data_out_386  (wire_weight_from_rom[386]),
			.data_out_387  (wire_weight_from_rom[387]),
			.data_out_388  (wire_weight_from_rom[388]),
			.data_out_389  (wire_weight_from_rom[389]),
			.data_out_390  (wire_weight_from_rom[390]),
			.data_out_391  (wire_weight_from_rom[391]),
			.data_out_392  (wire_weight_from_rom[392]),
			.data_out_393  (wire_weight_from_rom[393]),
			.data_out_394  (wire_weight_from_rom[394]),
			.data_out_395  (wire_weight_from_rom[395]),
			.data_out_396  (wire_weight_from_rom[396]),
			.data_out_397  (wire_weight_from_rom[397]),
			.data_out_398  (wire_weight_from_rom[398]),
			.data_out_399  (wire_weight_from_rom[399]),
			.data_out_400  (wire_weight_from_rom[400]),
			.data_out_401  (wire_weight_from_rom[401]),
			.data_out_402  (wire_weight_from_rom[402]),
			.data_out_403  (wire_weight_from_rom[403]),
			.data_out_404  (wire_weight_from_rom[404]),
			.data_out_405  (wire_weight_from_rom[405]),
			.data_out_406  (wire_weight_from_rom[406]),
			.data_out_407  (wire_weight_from_rom[407]),
			.data_out_408  (wire_weight_from_rom[408]),
			.data_out_409  (wire_weight_from_rom[409]),
			.data_out_410  (wire_weight_from_rom[410]),
			.data_out_411  (wire_weight_from_rom[411]),
			.data_out_412  (wire_weight_from_rom[412]),
			.data_out_413  (wire_weight_from_rom[413]),
			.data_out_414  (wire_weight_from_rom[414]),
			.data_out_415  (wire_weight_from_rom[415]),
			.data_out_416  (wire_weight_from_rom[416]),
			.data_out_417  (wire_weight_from_rom[417]),
			.data_out_418  (wire_weight_from_rom[418]),
			.data_out_419  (wire_weight_from_rom[419]),
			.data_out_420  (wire_weight_from_rom[420]),
			.data_out_421  (wire_weight_from_rom[421]),
			.data_out_422  (wire_weight_from_rom[422]),
			.data_out_423  (wire_weight_from_rom[423]),
			.data_out_424  (wire_weight_from_rom[424]),
			.data_out_425  (wire_weight_from_rom[425]),
			.data_out_426  (wire_weight_from_rom[426]),
			.data_out_427  (wire_weight_from_rom[427]),
			.data_out_428  (wire_weight_from_rom[428]),
			.data_out_429  (wire_weight_from_rom[429]),
			.data_out_430  (wire_weight_from_rom[430]),
			.data_out_431  (wire_weight_from_rom[431]),
			.data_out_432  (wire_weight_from_rom[432]),
			.data_out_433  (wire_weight_from_rom[433]),
			.data_out_434  (wire_weight_from_rom[434]),
			.data_out_435  (wire_weight_from_rom[435]),
			.data_out_436  (wire_weight_from_rom[436]),
			.data_out_437  (wire_weight_from_rom[437]),
			.data_out_438  (wire_weight_from_rom[438]),
			.data_out_439  (wire_weight_from_rom[439]),
			.data_out_440  (wire_weight_from_rom[440]),
			.data_out_441  (wire_weight_from_rom[441]),
			.data_out_442  (wire_weight_from_rom[442]),
			.data_out_443  (wire_weight_from_rom[443]),
			.data_out_444  (wire_weight_from_rom[444]),
			.data_out_445  (wire_weight_from_rom[445]),
			.data_out_446  (wire_weight_from_rom[446]),
			.data_out_447  (wire_weight_from_rom[447]),
			.data_out_448  (wire_weight_from_rom[448]),
			.data_out_449  (wire_weight_from_rom[449]),
			.data_out_450  (wire_weight_from_rom[450]),
			.data_out_451  (wire_weight_from_rom[451]),
			.data_out_452  (wire_weight_from_rom[452]),
			.data_out_453  (wire_weight_from_rom[453]),
			.data_out_454  (wire_weight_from_rom[454]),
			.data_out_455  (wire_weight_from_rom[455]),
			.data_out_456  (wire_weight_from_rom[456]),
			.data_out_457  (wire_weight_from_rom[457]),
			.data_out_458  (wire_weight_from_rom[458]),
			.data_out_459  (wire_weight_from_rom[459]),
			.data_out_460  (wire_weight_from_rom[460]),
			.data_out_461  (wire_weight_from_rom[461]),
			.data_out_462  (wire_weight_from_rom[462]),
			.data_out_463  (wire_weight_from_rom[463]),
			.data_out_464  (wire_weight_from_rom[464]),
			.data_out_465  (wire_weight_from_rom[465]),
			.data_out_466  (wire_weight_from_rom[466]),
			.data_out_467  (wire_weight_from_rom[467]),
			.data_out_468  (wire_weight_from_rom[468]),
			.data_out_469  (wire_weight_from_rom[469]),
			.data_out_470  (wire_weight_from_rom[470]),
			.data_out_471  (wire_weight_from_rom[471]),
			.data_out_472  (wire_weight_from_rom[472]),
			.data_out_473  (wire_weight_from_rom[473]),
			.data_out_474  (wire_weight_from_rom[474]),
			.data_out_475  (wire_weight_from_rom[475]),
			.data_out_476  (wire_weight_from_rom[476]),
			.data_out_477  (wire_weight_from_rom[477]),
			.data_out_478  (wire_weight_from_rom[478]),
			.data_out_479  (wire_weight_from_rom[479]),
			.data_out_480  (wire_weight_from_rom[480]),
			.data_out_481  (wire_weight_from_rom[481]),
			.data_out_482  (wire_weight_from_rom[482]),
			.data_out_483  (wire_weight_from_rom[483]),
			.data_out_484  (wire_weight_from_rom[484]),
			.data_out_485  (wire_weight_from_rom[485]),
			.data_out_486  (wire_weight_from_rom[486]),
			.data_out_487  (wire_weight_from_rom[487]),
			.data_out_488  (wire_weight_from_rom[488]),
			.data_out_489  (wire_weight_from_rom[489]),
			.data_out_490  (wire_weight_from_rom[490]),
			.data_out_491  (wire_weight_from_rom[491]),
			.data_out_492  (wire_weight_from_rom[492]),
			.data_out_493  (wire_weight_from_rom[493]),
			.data_out_494  (wire_weight_from_rom[494]),
			.data_out_495  (wire_weight_from_rom[495]),
			.data_out_496  (wire_weight_from_rom[496]),
			.data_out_497  (wire_weight_from_rom[497]),
			.data_out_498  (wire_weight_from_rom[498]),
			.data_out_499  (wire_weight_from_rom[499]),
			.data_out_500  (wire_weight_from_rom[500]),
			.data_out_501  (wire_weight_from_rom[501]),
			.data_out_502  (wire_weight_from_rom[502]),
			.data_out_503  (wire_weight_from_rom[503]),
			.data_out_504  (wire_weight_from_rom[504]),
			.data_out_505  (wire_weight_from_rom[505]),
			.data_out_506  (wire_weight_from_rom[506]),
			.data_out_507  (wire_weight_from_rom[507]),
			.data_out_508  (wire_weight_from_rom[508]),
			.data_out_509  (wire_weight_from_rom[509]),
			.data_out_510  (wire_weight_from_rom[510]),
			.data_out_511  (wire_weight_from_rom[511]),
			.data_out_512  (wire_weight_from_rom[512]),
			.data_out_513  (wire_weight_from_rom[513]),
			.data_out_514  (wire_weight_from_rom[514]),
			.data_out_515  (wire_weight_from_rom[515]),
			.data_out_516  (wire_weight_from_rom[516]),
			.data_out_517  (wire_weight_from_rom[517]),
			.data_out_518  (wire_weight_from_rom[518]),
			.data_out_519  (wire_weight_from_rom[519]),
			.data_out_520  (wire_weight_from_rom[520]),
			.data_out_521  (wire_weight_from_rom[521]),
			.data_out_522  (wire_weight_from_rom[522]),
			.data_out_523  (wire_weight_from_rom[523]),
			.data_out_524  (wire_weight_from_rom[524]),
			.data_out_525  (wire_weight_from_rom[525]),
			.data_out_526  (wire_weight_from_rom[526]),
			.data_out_527  (wire_weight_from_rom[527]),
			.data_out_528  (wire_weight_from_rom[528]),
			.data_out_529  (wire_weight_from_rom[529]),
			.data_out_530  (wire_weight_from_rom[530]),
			.data_out_531  (wire_weight_from_rom[531]),
			.data_out_532  (wire_weight_from_rom[532]),
			.data_out_533  (wire_weight_from_rom[533]),
			.data_out_534  (wire_weight_from_rom[534]),
			.data_out_535  (wire_weight_from_rom[535]),
			.data_out_536  (wire_weight_from_rom[536]),
			.data_out_537  (wire_weight_from_rom[537]),
			.data_out_538  (wire_weight_from_rom[538]),
			.data_out_539  (wire_weight_from_rom[539]),
			.data_out_540  (wire_weight_from_rom[540]),
			.data_out_541  (wire_weight_from_rom[541]),
			.data_out_542  (wire_weight_from_rom[542]),
			.data_out_543  (wire_weight_from_rom[543]),
			.data_out_544  (wire_weight_from_rom[544]),
			.data_out_545  (wire_weight_from_rom[545]),
			.data_out_546  (wire_weight_from_rom[546]),
			.data_out_547  (wire_weight_from_rom[547]),
			.data_out_548  (wire_weight_from_rom[548]),
			.data_out_549  (wire_weight_from_rom[549]),
			.data_out_550  (wire_weight_from_rom[550]),
			.data_out_551  (wire_weight_from_rom[551]),
			.data_out_552  (wire_weight_from_rom[552]),
			.data_out_553  (wire_weight_from_rom[553]),
			.data_out_554  (wire_weight_from_rom[554]),
			.data_out_555  (wire_weight_from_rom[555]),
			.data_out_556  (wire_weight_from_rom[556]),
			.data_out_557  (wire_weight_from_rom[557]),
			.data_out_558  (wire_weight_from_rom[558]),
			.data_out_559  (wire_weight_from_rom[559]),
			.data_out_560  (wire_weight_from_rom[560]),
			.data_out_561  (wire_weight_from_rom[561]),
			.data_out_562  (wire_weight_from_rom[562]),
			.data_out_563  (wire_weight_from_rom[563]),
			.data_out_564  (wire_weight_from_rom[564]),
			.data_out_565  (wire_weight_from_rom[565]),
			.data_out_566  (wire_weight_from_rom[566]),
			.data_out_567  (wire_weight_from_rom[567]),
			.data_out_568  (wire_weight_from_rom[568]),
			.data_out_569  (wire_weight_from_rom[569]),
			.data_out_570  (wire_weight_from_rom[570]),
			.data_out_571  (wire_weight_from_rom[571]),
			.data_out_572  (wire_weight_from_rom[572]),
			.data_out_573  (wire_weight_from_rom[573]),
			.data_out_574  (wire_weight_from_rom[574]),
			.data_out_575  (wire_weight_from_rom[575]),
			.data_out_576  (wire_weight_from_rom[576]),
			.data_out_577  (wire_weight_from_rom[577]),
			.data_out_578  (wire_weight_from_rom[578]),
			.data_out_579  (wire_weight_from_rom[579]),
			.data_out_580  (wire_weight_from_rom[580]),
			.data_out_581  (wire_weight_from_rom[581]),
			.data_out_582  (wire_weight_from_rom[582]),
			.data_out_583  (wire_weight_from_rom[583]),
			.data_out_584  (wire_weight_from_rom[584]),
			.data_out_585  (wire_weight_from_rom[585]),
			.data_out_586  (wire_weight_from_rom[586]),
			.data_out_587  (wire_weight_from_rom[587]),
			.data_out_588  (wire_weight_from_rom[588]),
			.data_out_589  (wire_weight_from_rom[589]),
			.data_out_590  (wire_weight_from_rom[590]),
			.data_out_591  (wire_weight_from_rom[591]),
			.data_out_592  (wire_weight_from_rom[592]),
			.data_out_593  (wire_weight_from_rom[593]),
			.data_out_594  (wire_weight_from_rom[594]),
			.data_out_595  (wire_weight_from_rom[595]),
			.data_out_596  (wire_weight_from_rom[596]),
			.data_out_597  (wire_weight_from_rom[597]),
			.data_out_598  (wire_weight_from_rom[598]),
			.data_out_599  (wire_weight_from_rom[599]),
			.data_out_600  (wire_weight_from_rom[600]),
			.data_out_601  (wire_weight_from_rom[601]),
			.data_out_602  (wire_weight_from_rom[602]),
			.data_out_603  (wire_weight_from_rom[603]),
			.data_out_604  (wire_weight_from_rom[604]),
			.data_out_605  (wire_weight_from_rom[605]),
			.data_out_606  (wire_weight_from_rom[606]),
			.data_out_607  (wire_weight_from_rom[607]),
			.data_out_608  (wire_weight_from_rom[608]),
			.data_out_609  (wire_weight_from_rom[609]),
			.data_out_610  (wire_weight_from_rom[610]),
			.data_out_611  (wire_weight_from_rom[611]),
			.data_out_612  (wire_weight_from_rom[612]),
			.data_out_613  (wire_weight_from_rom[613]),
			.data_out_614  (wire_weight_from_rom[614]),
			.data_out_615  (wire_weight_from_rom[615]),
			.data_out_616  (wire_weight_from_rom[616]),
			.data_out_617  (wire_weight_from_rom[617]),
			.data_out_618  (wire_weight_from_rom[618]),
			.data_out_619  (wire_weight_from_rom[619]),
			.data_out_620  (wire_weight_from_rom[620]),
			.data_out_621  (wire_weight_from_rom[621]),
			.data_out_622  (wire_weight_from_rom[622]),
			.data_out_623  (wire_weight_from_rom[623]),
			.data_out_624  (wire_weight_from_rom[624]),
			.data_out_625  (wire_weight_from_rom[625]),
			.data_out_626  (wire_weight_from_rom[626]),
			.data_out_627  (wire_weight_from_rom[627]),
			.data_out_628  (wire_weight_from_rom[628]),
			.data_out_629  (wire_weight_from_rom[629]),
			.data_out_630  (wire_weight_from_rom[630]),
			.data_out_631  (wire_weight_from_rom[631]),
			.data_out_632  (wire_weight_from_rom[632]),
			.data_out_633  (wire_weight_from_rom[633]),
			.data_out_634  (wire_weight_from_rom[634]),
			.data_out_635  (wire_weight_from_rom[635]),
			.data_out_636  (wire_weight_from_rom[636]),
			.data_out_637  (wire_weight_from_rom[637]),
			.data_out_638  (wire_weight_from_rom[638]),
			.data_out_639  (wire_weight_from_rom[639]),
			.data_out_640  (wire_weight_from_rom[640]),
			.data_out_641  (wire_weight_from_rom[641]),
			.data_out_642  (wire_weight_from_rom[642]),
			.data_out_643  (wire_weight_from_rom[643]),
			.data_out_644  (wire_weight_from_rom[644]),
			.data_out_645  (wire_weight_from_rom[645]),
			.data_out_646  (wire_weight_from_rom[646]),
			.data_out_647  (wire_weight_from_rom[647]),
			.data_out_648  (wire_weight_from_rom[648]),
			.data_out_649  (wire_weight_from_rom[649]),
			.data_out_650  (wire_weight_from_rom[650]),
			.data_out_651  (wire_weight_from_rom[651]),
			.data_out_652  (wire_weight_from_rom[652]),
			.data_out_653  (wire_weight_from_rom[653]),
			.data_out_654  (wire_weight_from_rom[654]),
			.data_out_655  (wire_weight_from_rom[655]),
			.data_out_656  (wire_weight_from_rom[656]),
			.data_out_657  (wire_weight_from_rom[657]),
			.data_out_658  (wire_weight_from_rom[658]),
			.data_out_659  (wire_weight_from_rom[659]),
			.data_out_660  (wire_weight_from_rom[660]),
			.data_out_661  (wire_weight_from_rom[661]),
			.data_out_662  (wire_weight_from_rom[662]),
			.data_out_663  (wire_weight_from_rom[663]),
			.data_out_664  (wire_weight_from_rom[664]),
			.data_out_665  (wire_weight_from_rom[665]),
			.data_out_666  (wire_weight_from_rom[666]),
			.data_out_667  (wire_weight_from_rom[667]),
			.data_out_668  (wire_weight_from_rom[668]),
			.data_out_669  (wire_weight_from_rom[669]),
			.data_out_670  (wire_weight_from_rom[670]),
			.data_out_671  (wire_weight_from_rom[671]),
			.data_out_672  (wire_weight_from_rom[672]),
			.data_out_673  (wire_weight_from_rom[673]),
			.data_out_674  (wire_weight_from_rom[674]),
			.data_out_675  (wire_weight_from_rom[675]),
			.data_out_676  (wire_weight_from_rom[676]),
			.data_out_677  (wire_weight_from_rom[677]),
			.data_out_678  (wire_weight_from_rom[678]),
			.data_out_679  (wire_weight_from_rom[679]),
			.data_out_680  (wire_weight_from_rom[680]),
			.data_out_681  (wire_weight_from_rom[681]),
			.data_out_682  (wire_weight_from_rom[682]),
			.data_out_683  (wire_weight_from_rom[683]),
			.data_out_684  (wire_weight_from_rom[684]),
			.data_out_685  (wire_weight_from_rom[685]),
			.data_out_686  (wire_weight_from_rom[686]),
			.data_out_687  (wire_weight_from_rom[687]),
			.data_out_688  (wire_weight_from_rom[688]),
			.data_out_689  (wire_weight_from_rom[689]),
			.data_out_690  (wire_weight_from_rom[690]),
			.data_out_691  (wire_weight_from_rom[691]),
			.data_out_692  (wire_weight_from_rom[692]),
			.data_out_693  (wire_weight_from_rom[693]),
			.data_out_694  (wire_weight_from_rom[694]),
			.data_out_695  (wire_weight_from_rom[695]),
			.data_out_696  (wire_weight_from_rom[696]),
			.data_out_697  (wire_weight_from_rom[697]),
			.data_out_698  (wire_weight_from_rom[698]),
			.data_out_699  (wire_weight_from_rom[699]),
			.data_out_700  (wire_weight_from_rom[700]),
			.data_out_701  (wire_weight_from_rom[701]),
			.data_out_702  (wire_weight_from_rom[702]),
			.data_out_703  (wire_weight_from_rom[703]),
			.data_out_704  (wire_weight_from_rom[704]),
			.data_out_705  (wire_weight_from_rom[705]),
			.data_out_706  (wire_weight_from_rom[706]),
			.data_out_707  (wire_weight_from_rom[707]),
			.data_out_708  (wire_weight_from_rom[708]),
			.data_out_709  (wire_weight_from_rom[709]),
			.data_out_710  (wire_weight_from_rom[710]),
			.data_out_711  (wire_weight_from_rom[711]),
			.data_out_712  (wire_weight_from_rom[712]),
			.data_out_713  (wire_weight_from_rom[713]),
			.data_out_714  (wire_weight_from_rom[714]),
			.data_out_715  (wire_weight_from_rom[715]),
			.data_out_716  (wire_weight_from_rom[716]),
			.data_out_717  (wire_weight_from_rom[717]),
			.data_out_718  (wire_weight_from_rom[718]),
			.data_out_719  (wire_weight_from_rom[719]),
			.data_out_720  (wire_weight_from_rom[720]),
			.data_out_721  (wire_weight_from_rom[721]),
			.data_out_722  (wire_weight_from_rom[722]),
			.data_out_723  (wire_weight_from_rom[723]),
			.data_out_724  (wire_weight_from_rom[724]),
			.data_out_725  (wire_weight_from_rom[725]),
			.data_out_726  (wire_weight_from_rom[726]),
			.data_out_727  (wire_weight_from_rom[727]),
			.data_out_728  (wire_weight_from_rom[728]),
			.data_out_729  (wire_weight_from_rom[729]),
			.data_out_730  (wire_weight_from_rom[730]),
			.data_out_731  (wire_weight_from_rom[731]),
			.data_out_732  (wire_weight_from_rom[732]),
			.data_out_733  (wire_weight_from_rom[733]),
			.data_out_734  (wire_weight_from_rom[734]),
			.data_out_735  (wire_weight_from_rom[735]),
			.data_out_736  (wire_weight_from_rom[736]),
			.data_out_737  (wire_weight_from_rom[737]),
			.data_out_738  (wire_weight_from_rom[738]),
			.data_out_739  (wire_weight_from_rom[739])

		
		
		
	);
	
	
	
	// ======================== HIDDEN LAYER START ===============================
	
	genvar ii;
	generate
		for (ii = 0; ii < 10; ii = ii + 1) begin : gen_hidden_layer
			NPU_dotproduct hidden_layer_neuron(
			.clk(clk),
			.reset(reset),
			.data(data_in),
			.wire_weight_from_rom_63  (wire_weight_from_rom[(ii*64) + 0 ]     ),
			.wire_weight_from_rom_62  (wire_weight_from_rom[(ii*64) + 1 ]     ),
			.wire_weight_from_rom_61  (wire_weight_from_rom[(ii*64) + 2 ]     ),
			.wire_weight_from_rom_60  (wire_weight_from_rom[(ii*64) + 3 ]     ),
			.wire_weight_from_rom_59  (wire_weight_from_rom[(ii*64) + 4 ]     ),
			.wire_weight_from_rom_58  (wire_weight_from_rom[(ii*64) + 5 ]     ),
			.wire_weight_from_rom_57  (wire_weight_from_rom[(ii*64) + 6 ]     ),
			.wire_weight_from_rom_56  (wire_weight_from_rom[(ii*64) + 7 ]     ),
			.wire_weight_from_rom_55  (wire_weight_from_rom[(ii*64) + 8 ]     ),
			.wire_weight_from_rom_54  (wire_weight_from_rom[(ii*64) + 9 ]     ),
			.wire_weight_from_rom_53  (wire_weight_from_rom[(ii*64) + 10]     ),
			.wire_weight_from_rom_52  (wire_weight_from_rom[(ii*64) + 11]     ),
			.wire_weight_from_rom_51  (wire_weight_from_rom[(ii*64) + 12]     ),
			.wire_weight_from_rom_50  (wire_weight_from_rom[(ii*64) + 13]     ),
			.wire_weight_from_rom_49  (wire_weight_from_rom[(ii*64) + 14]     ),
			.wire_weight_from_rom_48  (wire_weight_from_rom[(ii*64) + 15]     ),
			.wire_weight_from_rom_47  (wire_weight_from_rom[(ii*64) + 16]     ),
			.wire_weight_from_rom_46  (wire_weight_from_rom[(ii*64) + 17]     ),
			.wire_weight_from_rom_45  (wire_weight_from_rom[(ii*64) + 18]     ),
			.wire_weight_from_rom_44  (wire_weight_from_rom[(ii*64) + 19]     ),
			.wire_weight_from_rom_43  (wire_weight_from_rom[(ii*64) + 20]     ),
			.wire_weight_from_rom_42  (wire_weight_from_rom[(ii*64) + 21]     ),
			.wire_weight_from_rom_41  (wire_weight_from_rom[(ii*64) + 22]     ),
			.wire_weight_from_rom_40  (wire_weight_from_rom[(ii*64) + 23]     ),
			.wire_weight_from_rom_39  (wire_weight_from_rom[(ii*64) + 24]     ),
			.wire_weight_from_rom_38  (wire_weight_from_rom[(ii*64) + 25]     ),
			.wire_weight_from_rom_37  (wire_weight_from_rom[(ii*64) + 26]     ),
			.wire_weight_from_rom_36  (wire_weight_from_rom[(ii*64) + 27]     ),
			.wire_weight_from_rom_35  (wire_weight_from_rom[(ii*64) + 28]     ),
			.wire_weight_from_rom_34  (wire_weight_from_rom[(ii*64) + 29]     ),
			.wire_weight_from_rom_33  (wire_weight_from_rom[(ii*64) + 30]     ),
			.wire_weight_from_rom_32  (wire_weight_from_rom[(ii*64) + 31]     ),
			.wire_weight_from_rom_31  (wire_weight_from_rom[(ii*64) + 32]     ),
			.wire_weight_from_rom_30  (wire_weight_from_rom[(ii*64) + 33]     ),
			.wire_weight_from_rom_29  (wire_weight_from_rom[(ii*64) + 34]     ),
			.wire_weight_from_rom_28  (wire_weight_from_rom[(ii*64) + 35]     ),
			.wire_weight_from_rom_27  (wire_weight_from_rom[(ii*64) + 36]     ),
			.wire_weight_from_rom_26  (wire_weight_from_rom[(ii*64) + 37]     ),
			.wire_weight_from_rom_25  (wire_weight_from_rom[(ii*64) + 38]     ),
			.wire_weight_from_rom_24  (wire_weight_from_rom[(ii*64) + 39]     ),
			.wire_weight_from_rom_23  (wire_weight_from_rom[(ii*64) + 40]     ),
			.wire_weight_from_rom_22  (wire_weight_from_rom[(ii*64) + 41]     ),
			.wire_weight_from_rom_21  (wire_weight_from_rom[(ii*64) + 42]     ),
			.wire_weight_from_rom_20  (wire_weight_from_rom[(ii*64) + 43]     ),
			.wire_weight_from_rom_19  (wire_weight_from_rom[(ii*64) + 44]     ),
			.wire_weight_from_rom_18  (wire_weight_from_rom[(ii*64) + 45]     ),
			.wire_weight_from_rom_17  (wire_weight_from_rom[(ii*64) + 46]     ),
			.wire_weight_from_rom_16  (wire_weight_from_rom[(ii*64) + 47]     ),
			.wire_weight_from_rom_15  (wire_weight_from_rom[(ii*64) + 48]     ),
			.wire_weight_from_rom_14  (wire_weight_from_rom[(ii*64) + 49]     ),
			.wire_weight_from_rom_13  (wire_weight_from_rom[(ii*64) + 50]     ),
			.wire_weight_from_rom_12  (wire_weight_from_rom[(ii*64) + 51]     ),
			.wire_weight_from_rom_11  (wire_weight_from_rom[(ii*64) + 52]     ),
			.wire_weight_from_rom_10  (wire_weight_from_rom[(ii*64) + 53]     ),
			.wire_weight_from_rom_9   (wire_weight_from_rom[(ii*64) + 54]     ),
			.wire_weight_from_rom_8   (wire_weight_from_rom[(ii*64) + 55]     ),
			.wire_weight_from_rom_7   (wire_weight_from_rom[(ii*64) + 56]     ),
			.wire_weight_from_rom_6   (wire_weight_from_rom[(ii*64) + 57]     ),
			.wire_weight_from_rom_5   (wire_weight_from_rom[(ii*64) + 58]     ),
			.wire_weight_from_rom_4   (wire_weight_from_rom[(ii*64) + 59]     ),
			.wire_weight_from_rom_3   (wire_weight_from_rom[(ii*64) + 60]     ),
			.wire_weight_from_rom_2   (wire_weight_from_rom[(ii*64) + 61]     ),
			.wire_weight_from_rom_1   (wire_weight_from_rom[(ii*64) + 62]     ),
			.wire_weight_from_rom_0   (wire_weight_from_rom[(ii*64) + 63]     ),
			
			.result(wire_hiddenlayer_neuron_result[ii])
			
		);
		end
	endgenerate

	
	
	// Activation Function: ReLu
	genvar j;
	generate
		for (j = 0 ; j<10 ; j = j+1) begin: gen_ReLu
			ReLu ReLu (
				.data_in(wire_hiddenlayer_neuron_result[j]),
				.result(wire_ReLu_result[j])
			);
		end
	endgenerate
	
	// ======================== HIDDEN LAYER END ===============================




	// ======================== OUTPUT LAYER START ===============================
	
	genvar i;
	generate
		for (i = 0; i < 10; i = i + 1) begin: output_neuron
			Output_Layer_Neuron Output_Layer_Neuron(
			.clk    (clk), 
			.reset  (reset),
			.ReLu0  (wire_ReLu_result[0]),
			.ReLu1  (wire_ReLu_result[1]),
			.ReLu2  (wire_ReLu_result[2]),
			.ReLu3  (wire_ReLu_result[3]),
			.ReLu4  (wire_ReLu_result[4]),
			.ReLu5  (wire_ReLu_result[5]),
			.ReLu6  (wire_ReLu_result[6]),
			.ReLu7  (wire_ReLu_result[7]),
			.ReLu8  (wire_ReLu_result[8]),
			.ReLu9  (wire_ReLu_result[9]),
			
			
			
			.Weight0(wire_weight_from_rom[(i*10)+640]),
			.Weight1(wire_weight_from_rom[(i*10)+641]),
			.Weight2(wire_weight_from_rom[(i*10)+642]),
			.Weight3(wire_weight_from_rom[(i*10)+643]),
			.Weight4(wire_weight_from_rom[(i*10)+644]),
			.Weight5(wire_weight_from_rom[(i*10)+645]),
			.Weight6(wire_weight_from_rom[(i*10)+646]),
			.Weight7(wire_weight_from_rom[(i*10)+647]),
			.Weight8(wire_weight_from_rom[(i*10)+648]),
			.Weight9(wire_weight_from_rom[(i*10)+649]),
			

			.result (output_layer_neuron[i])
		);
		end
	endgenerate
		
		
		
		
		

	
	
	
	
	
	
	
	
	// ======================== OUTPUT LAYER END===============================
	
	
	// ======================== COMPARATOR START ===============================
	Max_Find_10_Bfloat16 Final_Inference(
		.input_0(output_layer_neuron[0]),
		.input_1(output_layer_neuron[1]),
		.input_2(output_layer_neuron[2]),
		.input_3(output_layer_neuron[3]),
		.input_4(output_layer_neuron[4]),
		.input_5(output_layer_neuron[5]),
		.input_6(output_layer_neuron[6]),
		.input_7(output_layer_neuron[7]),
		.input_8(output_layer_neuron[8]),
		.input_9(output_layer_neuron[9]),
		
		.result(final_inference)
	
	);
	
	
	
	// ======================== COMPARATOR END ===============================
	



   
endmodule
